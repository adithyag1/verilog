module fullpractb;
    reg a,b,c;
    wire S,C;

    fullprac uut(
        .a(a),
        .b(b),
        .c(c),
        .S(S),
        .C(C)
    )

    integer i,j,k;
    
endmodule 
    